library verilog;
use verilog.vl_types.all;
entity multiTest is
end multiTest;
