module DecryptionMonPro(n,d,c,clk,m);
					

input [31:0] n; //product of prime numbers
input [31:0] d; //private key
input [31:0] c; //cipher text
input clk;


output [31:0] m; //plain text
 
//instatiate all of the lower level modules here

endmodule
